module adder (input A, input  B, wire Q);


assign Q = A + B;


    
endmodule
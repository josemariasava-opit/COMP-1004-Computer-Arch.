module and_gate(input A, input B, output Q);

    assign Y = A & B;

endmodule